// Defines for ECP5 evaluation board
// `define SPI_FLASH
